��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CLogicOut�� 	 CTerminal   ��               �            x$�           ��    �
�  `(u)     	          �            t �0           ��    ��  CNAND
�  �x�y              @          
�  ����              @          
�  ����               �            �t��           ��    �
�  � �!              @          
�  �0�1              @          
�  ())     	          �            �4           ��    �
�  Pxey               �          
�  P�e�              @          
�  |���              @            dt|�           ��    �
�  �p�q              @          
�  ����              @          
�  x)y               �            �l�           ��    �
�  �p�q              @          
�  ����               �          
�  �x�y              @            �l��            ��    �
�  � pq              @          
�  � ��              @          
�  x1y     
          �            l�     $      ��    �
�  8pMq     
          �          
�  8�M�     
          �          
�  dxyy              @            Lld�     (      ��    �
�  � �!               �          
�  �0�1               �          
�  �(�)              @            ��4     ,      ��    �
�  ` �u �              @          
�  ` �u �              @          
�  � �� �               �            t �� �     0      ��    ��  CLogicIn�� 	 CLatchKey   � �     4   
�  $ �9 �              @             �$ �     7   ����     3�5�   I W     8   
�  $ P9 Q              @             L$ T     :   ����     �
�  (� =�               @          
�  (� =�               @          
�  T� i�                �            <� T�      <      ��    �
�  � � � �                �          
�  � � � �               @          
�  � � 	�               @            � � � �      @      ��    �
�  p � � �               @          
�  p � � �               @          
�  � � � �                �            � � � �      D      ��    3�5�   �   �      G   
�  , � A �               @            $ � , �      I   ����                   ���  CWire  ���      K�  ((a)     	 K�  ����       K�  ����      K�  �x�y      K�  �x��       K�  P�Q�       K�  ��Q�      K��� 
 CCrossOver  �t�|        �(��       K�  �(�)      K�U�  �t�|        �x�y      K�  �(�)      K�  �(�1       K�  � �)       K�  (xQy      K�  �x��       K�  �p�y       K�  ����       K�  � ���      K�U�  � |� �      U�  � l� t      U�  � L� T      U�  � � $        � � � �       K�  � � � �       K�U�  � |� �      U�  � |� �        h �� �      K�U�  � l� t      U�  f ll t      U�  � l� t        H p� q      K�U�  � L� T      U�  � L� T        h P� Q      K�U�  � � $        � � � Q       K�U�  � � $      U�  fl$      U�  � � $        �  �!      K�  � � � �       K�  xx�y      K�  �p�y       K�U�  f ll t        h Pi �       K�  8 Pi Q      K�U�  � |� �      U�  � l� t      U�  � L� T        �  � �       K�  H pI �       K�  8 �I �      K�  H �a �      K�  0p1y      
 K�  0p9q     
 K�  0x1�      
 K�  0�9�     
 K�  h0�1      K�U�  fl$        h� i1       K�  ` �a �       K�  ` �a �       K�  (� )�        K�  (� )�        K�  � )�       K�  p � q �        K�  p � q �        K�  @ � q �                     �                             L   M   P   N    L  \   [    M  ]   R    Q  _   ^    ]   z   ! ` ! " " X $ k $ % h % & & � ( � ( ) � ) * * y , t , - � - . . W 0 � 0 1 � 1 2 2 ~ 7 7 � : : } < � < = � = > > � @ x @ A r A B B � D � D E � E F F g I I �     O   N Q  P O  S T R T Y Z S . T X V " ^ W \ Z   [   _   X ! a b ` b i b l b p b u x a F b h c h  { % k d k | k � � $ o e o � } r r w A o t f t � t s ~ , g @ * z   y { m o h : { ~ j ~ n ~ q t 2 k � 7 � � � � � � ( & � � ) � - � v > � � 1 0 � < � � = B � � E D � I �             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 