��  CCircuit��  CSerializeHack           ��  CPart              ���  CNAND�� 	 CTerminal  h�}�               �          
�  h�}�               �          
�  ����              @            |���           ��    �� 	 CLogicOut
�  ����               �            ����           ��    �
�  �H�I               �            �@�P           ��    ��  CLogicIn�� 	 CLatchKey  H�X�        
�  d�y�              @            \�d�        ����     ��  HQX_        
�  dXyY              @            \Td\        ����     ��  P`        
�  l�	              @            dl        ����     �
�  ���              @          
�  ���              @          
�  $�9�               �            �$�           ��    �
�  ���     
          �          
�  ���              @          
�  �1�              @            |�     #      ��    �
�  �@�A              @          
�  �P�Q              @          
�  H)I               �            �<T     '      ��    �
�  � �     	         @          
�  ��               �          
�  !	              @            ��      +      ��    �
�  `puq              @          
�  `�u�              @          
�  �x�y               �            tl��     /      ��    �
�  X8m9     	         @          
�  XHmI     	         @          
�  �@�A               �            l4�L     3      ��    �
�  X m               �          
�  Xm               �          
�  ��	     	         @            l� �     7      ��    �
�  ����              @          
�  ����              @          
�  ���               �            ����     ;      ��    �
�  �p�q              @          
�  ����              @          
�  xy               �            �l�     ?      ��    �
�  �8�9     
          �          
�  �H�I              @          
�  @A              @            �4L     C      ��    �
�  � �              @          
�  ��              @          
�  	     
          �            ��      G      ��                  ���  CWire�� 
 CCrossOver  VD\L        (HiI      K�M�  VD\L      M�  V\\d        X Y�       K�M�  f\ld        hHi�       K�  h���      K�M�  f\ld      M�  �\�d      M�  V\\d        �`�a      K�  �@�A      K�  �@�a       K�  �H�a       K�  �x�y      K�M�  �\�d      M�  �� �        �� ��      
 K�  ����      K�  ����       K�  ����      K�  ����       K�  ��A�      K�  @�A�       K�  0�A�      K�  ����      K�  ����       K�  ����      K�  � 	      
 K�  � ��      
 K�  ����     
 K�M�  �� �        � �     	 K�  ��!       K�  �0�A       K�  �@�Q       K�  �P�Q      K�   1	      K�M�  .4$        011       K�  �011      K�M�  .4$        � Y!      K�  �@�A      K�  8�Y�      K�  ��      K�  � �	      	 K�  h�i�       K�  h�i�       K�  `�i�      K�  `�a�       K�  `�i�      K�  �x��       K�  h���      K�  x�y�       K�  x�Y�      K�M�  �l�t        �H��       K�  ��Q�      K�  X�Y�       K�  X�a�      K�  PpQ�       K�  �H�I      K�  xH�I      K�M�  �l�t        xp�q      K�  Ppaq      K�  HI�       K�M�  >|D�        @ A�       K�  P(Q9      	 K�  P8QI      	 K�  PHYI     	 K�  ��)      	 K�  P(�)     	 K�  P8Y9     	 K�  x�       K�M�  .|4�      M�  >|D�        �I�      K�M�  .|4�        0@1�       K�  HY      K�  �A�      K�  @ Y      K�  ����       K�  ����       K�  ����      K�  ����       K�  ����      K�  @1A      K�  ��1�      K�  ����      K�  �p�q      K�  �p��       K�  xpy�       K�  xHyY       K�  �8�9     
 K�  �(�9      
 K�  �()     
 K�  )      
 K�  ��	      K�  ��	      K�  ��       K�  ��      K�  � �	                     �                             }   �    g  T   [    �   �   �  `    b   ! ! z # l # $ i $ % % f ' y ' ( r ( ) ) L + m + , { , - - s / � / 0 � 0 1 1 \ 3 � 3 4 � 4 5 5 Y 7 � 7 8 � 8 9 9 � ; � ; < � < = = � ? � ? @ � @ A A � C � C D � D E E � G � G H � H I I � L P ) R O N O X w z R V L T R  U S U ^ U Q Z [ 5 Z Y U  U 1 � ] W ] n k l c  ` b a   d a c e f d % e  h i g h $ k I j ] ] # m _ | + { w v y p r q ( - t t x s v p t w u o O q ' ! O o , m 9 ~  �  � }  � �  \ � ~ �  � � � � � � � � � � � � 0 � � � D � � � � � � � / � � � � � � � � � � � 4 | � � � � 3 A � � � � � � � � � � � � 8 = � � 7 � ; � � � � � � � < E � � � � @ � ? � � � � �  � C � � � � j � � �  � � � � H G �             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 